library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;



package dadda_package is

	constant k: integer:=32;    --operand bits
	constant k_row:  integer:=33;	 --bits in the row k+1 bits
	--type array_level1 is array (0 to 16) of std_logic_vector(63 downto 0); -- matrix of layer 1
	


end package dadda_package;